netcdf tst_string_data {
dimensions:
	line = 5 ;
variables:
	string description(line) ;
		description:_FillValue = "" ;
data:

 description = "first string", "second string", "third string", _, 
    "last string" ;
}
