netcdf tst_opaque_data {
types:
  opaque(11) raw_obs_t ;
dimensions:
	time = 5 ;
variables:
	raw_obs_t raw_obs(time) ;
		raw_obs_t raw_obs:_FillValue = cafebabecafebabecafeba ;
data:

 raw_obs = 0102030405060708090a0b, aabbccddeeffeeddccbbaa, 
    ffffffffffffffffffffff, _, cf0defaced0cafe0facade ;
}
