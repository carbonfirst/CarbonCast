netcdf tst_solar_1 {
dimensions:
	length_of_name = 2 ;

// global attributes:
		:Number_of_vogons = 2dub, 23dub, 230dub ;
		:Number_of_vogon_poems = 23232244UL, 1214124123423UL, 2353424234UL ;

group: solar_system {

  group: Earth {

    // global attributes:
    		:alien_concept_number_which_cannot_be_understood_by_humans = -23232244L, 1214124123423L, -2353424234L ;

    group: Luna {
      variables:
      	int64 var_name(length_of_name) ;

      // global attributes:
      		:Vogon_Poem = "See, see the netCDF-filled sky\nMarvel at its big barf-green depths.\nTell me, Ed do you\nWonder why the yellow-bellied Snert ignores you?\nWhy its foobly stare\nmakes you feel ubiquitous obliquity.\nI can tell you, it is\nWorried by your HDF5-eating facial growth\nThat looks like\nA moldy pile of ASCII data.\nWhat\'s more, it knows\nYour redimensioning potting shed\nSmells of booger.\nEverything under the big netCDF-filled sky\nAsks why, why do you even bother?\nYou only charm software defects." ;
      data:

       var_name = 42, -42 ;
      } // group Luna
    } // group Earth
  } // group solar_system
}
